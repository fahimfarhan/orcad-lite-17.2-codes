CLANPER CKT 
VSIN a 0 SIN(0,10,1K, 0,0)
C1 A B 1
R1 B 0 1MEGA
VDC C 0 4
D1 C B DBREAK 
.MODEL DBREAK D
.PROBE
.TRAN 1U 4M
.END



