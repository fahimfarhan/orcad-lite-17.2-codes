TRANSIENT SIMULATION
* CMOS INVERTER
VIN 1 0 PULSE(0 5 0 1P 1P 5N 10N)
VDD 3 0 5
M2 2 1 3 3 PTYPE W=5U L= 2.5U
M1 2 1 0 0 NTYPE W = 5U L= 5U 

.MODEL PTYPE PMOS(KP=15U VTO=-1)
.MODEL NTYPE NMOS(KP=30U VTO=1) 

.PROBE
.TRAN 1N 20N 
.END

