MOSFET I-V CHARACTERISTICS
m1 1 2 0 0 ntype
.model ntype NMOS(VTO=1 kp=30u)
vgs 2 0 5
vds 1 0 5
.probe
.print dc i(vds)
.dc vds 0 5 0.5 vgs 0 5 1 
.end

